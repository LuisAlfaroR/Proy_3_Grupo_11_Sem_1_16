`timescale 1ns / 1ps

module font_rom
(
    input wire [10:0] addr,
	 input wire clk,
    output reg [23:0] data = 24'd0
);

//reg[23:0] data = 24'd0;

/*
always @(posedge clk) begin
	data_out <= data;
end
*/

always @ * begin
    data = 24'd0;
    case (addr)
      11'h0: data = 24'b000000000000000000000000;
      11'h1: data = 24'b000000000000000000000000;
      11'h2: data = 24'b000000000000000000000000;
      11'h3: data = 24'b000000000000000000000000;
      11'h4: data = 24'b000000000000000000000000;
      11'h5: data = 24'b000000000000000000000000;
      11'h6: data = 24'b000000000000000000000000;
      11'h7: data = 24'b000000000000000000000000;
      11'h8: data = 24'b000000000000000000000000;
      11'h9: data = 24'b111111111110000000000000;
      11'ha: data = 24'b111111111111100000000000;
      11'hb: data = 24'b111000000111110000000000;
      11'hc: data = 24'b111000000011111000000000;
      11'hd: data = 24'b111000000001111000000000;
      11'he: data = 24'b111000000000111000000000;
      11'hf: data = 24'b111000000000111100000000;
      11'h10: data = 24'b111000000000111100000000;
      11'h11: data = 24'b111000000000111100000000;
      11'h12: data = 24'b111000000000111100000000;
      11'h13: data = 24'b111000000000011100000000;
      11'h14: data = 24'b111000000000011100000000;
      11'h15: data = 24'b111000000000011100000000;
      11'h16: data = 24'b111000000000111100000000;
      11'h17: data = 24'b111000000000111100000000;
      11'h18: data = 24'b111000000000111100000000;
      11'h19: data = 24'b111000000000111100000000;
      11'h1a: data = 24'b111000000000111000000000;
      11'h1b: data = 24'b111000000001111000000000;
      11'h1c: data = 24'b111000000011110000000000;
      11'h1d: data = 24'b111000000111110000000000;
      11'h1e: data = 24'b111111111111100000000000;
      11'h1f: data = 24'b111111111110000000000000;
      11'h20: data = 24'b000000000000000000000000;
      11'h21: data = 24'b000000000000000000000000;
      11'h22: data = 24'b000000000000000000000000;
      11'h23: data = 24'b000000000000000000000000;
      11'h24: data = 24'b000000000000000000000000;
      11'h25: data = 24'b000000000000000000000000;
      11'h26: data = 24'b000000000000000000000000;
      11'h27: data = 24'b000000000000000000000000;
      11'h28: data = 24'b000000000000000000000000;
      11'h29: data = 24'b000000000000000000000000;
      11'h2a: data = 24'b000000000000000000000000;
      11'h2b: data = 24'b000000000000000000000000;
      11'h2c: data = 24'b000000000000000000000000;
      11'h2d: data = 24'b000000000000000000000000;
      11'h2e: data = 24'b000000000000000000000000;
      11'h2f: data = 24'b000000000000000000000000;

      11'h30: data = 24'b000000000000000000000000;
      11'h31: data = 24'b000000000000000000000000;
      11'h32: data = 24'b000000000000000000000000;
      11'h33: data = 24'b000000000000000000000000;
      11'h34: data = 24'b000000000000000000000000;
      11'h35: data = 24'b000000000000000000000000;
      11'h36: data = 24'b000000000000000000000000;
      11'h37: data = 24'b000000000000000000000000;
      11'h38: data = 24'b000000000000000000000000;
      11'h39: data = 24'b000000000000000000000000;
      11'h3a: data = 24'b000000000000000000000000;
      11'h3b: data = 24'b000000000000000000000000;
      11'h3c: data = 24'b000000111100000000000000;
      11'h3d: data = 24'b000000111100000000000000;
      11'h3e: data = 24'b000000000000000000000000;
      11'h3f: data = 24'b000000000000000000000000;
      11'h40: data = 24'b000000000000000000000000;
      11'h41: data = 24'b000000111100000000000000;
      11'h42: data = 24'b000000111100000000000000;
      11'h43: data = 24'b000000111100000000000000;
      11'h44: data = 24'b000000111100000000000000;
      11'h45: data = 24'b000000111100000000000000;
      11'h46: data = 24'b000000111100000000000000;
      11'h47: data = 24'b000000111100000000000000;
      11'h48: data = 24'b000000111100000000000000;
      11'h49: data = 24'b000000111100000000000000;
      11'h4a: data = 24'b000000111100000000000000;
      11'h4b: data = 24'b000000111100000000000000;
      11'h4c: data = 24'b000000111100000000000000;
      11'h4d: data = 24'b000000111100000000000000;
      11'h4e: data = 24'b000000111100000000000000;
      11'h4f: data = 24'b000000111100000000000000;
      11'h50: data = 24'b000000000000000000000000;
      11'h51: data = 24'b000000000000000000000000;
      11'h52: data = 24'b000000000000000000000000;
      11'h53: data = 24'b000000000000000000000000;
      11'h54: data = 24'b000000000000000000000000;
      11'h55: data = 24'b000000000000000000000000;
      11'h56: data = 24'b000000000000000000000000;
      11'h57: data = 24'b000000000000000000000000;
      11'h58: data = 24'b000000000000000000000000;
      11'h59: data = 24'b000000000000000000000000;
      11'h5a: data = 24'b000000000000000000000000;
      11'h5b: data = 24'b000000000000000000000000;
      11'h5c: data = 24'b000000000000000000000000;
      11'h5d: data = 24'b000000000000000000000000;
      11'h5e: data = 24'b000000000000000000000000;
      11'h5f: data = 24'b000000000000000000000000;

      11'h60: data = 24'b000000000000000000000000;
      11'h61: data = 24'b000000000000000000000000;
      11'h62: data = 24'b000000000000000000000000;
      11'h63: data = 24'b000000000000000000000000;
      11'h64: data = 24'b000000000000000000000000;
      11'h65: data = 24'b000000000000000000000000;
      11'h66: data = 24'b000000000000000000000000;
      11'h67: data = 24'b000000000000000000000000;
      11'h68: data = 24'b000000000000000000000000;
      11'h69: data = 24'b000000000000000000000000;
      11'h6a: data = 24'b000000000000000000000000;
      11'h6b: data = 24'b000000000000000000000000;
      11'h6c: data = 24'b000000000000000000000000;
      11'h6d: data = 24'b000000000000000000000000;
      11'h6e: data = 24'b000000000000000000000000;
      11'h6f: data = 24'b000011111111100000000000;
      11'h70: data = 24'b000111111111110000000000;
      11'h71: data = 24'b001111000011111000000000;
      11'h72: data = 24'b011110000001111000000000;
      11'h73: data = 24'b011110000001111000000000;
      11'h74: data = 24'b000000000001111000000000;
      11'h75: data = 24'b000000000011111000000000;
      11'h76: data = 24'b000011111111111000000000;
      11'h77: data = 24'b001111111111111000000000;
      11'h78: data = 24'b011111000001111000000000;
      11'h79: data = 24'b011110000001111000000000;
      11'h7a: data = 24'b111100000001111000000000;
      11'h7b: data = 24'b111100000001111000000000;
      11'h7c: data = 24'b011110000011111000000000;
      11'h7d: data = 24'b011110000111111000000000;
      11'h7e: data = 24'b001111111111111000000000;
      11'h7f: data = 24'b000111111100111100000000;
      11'h80: data = 24'b000000000000000000000000;
      11'h81: data = 24'b000000000000000000000000;
      11'h82: data = 24'b000000000000000000000000;
      11'h83: data = 24'b000000000000000000000000;
      11'h84: data = 24'b000000000000000000000000;
      11'h85: data = 24'b000000000000000000000000;
      11'h86: data = 24'b000000000000000000000000;
      11'h87: data = 24'b000000000000000000000000;
      11'h88: data = 24'b000000000000000000000000;
      11'h89: data = 24'b000000000000000000000000;
      11'h8a: data = 24'b000000000000000000000000;
      11'h8b: data = 24'b000000000000000000000000;
      11'h8c: data = 24'b000000000000000000000000;
      11'h8d: data = 24'b000000000000000000000000;
      11'h8e: data = 24'b000000000000000000000000;
      11'h8f: data = 24'b000000000000000000000000;

      11'h90: data = 24'b000000000000000000000000;
      11'h91: data = 24'b000000000000000000000000;
      11'h92: data = 24'b000000000000000000000000;
      11'h93: data = 24'b000000000000000000000000;
      11'h94: data = 24'b000000000000000000000000;
      11'h95: data = 24'b000000000000000000000000;
      11'h96: data = 24'b000000000000000000000000;
      11'h97: data = 24'b000000000000000000000000;
      11'h98: data = 24'b000000000000000000000000;
      11'h99: data = 24'b111100000001111000000000;
      11'h9a: data = 24'b111100000001111000000000;
      11'h9b: data = 24'b111100000001111000000000;
      11'h9c: data = 24'b111110000001111000000000;
      11'h9d: data = 24'b111110000011111000000000;
      11'h9e: data = 24'b111110000011111000000000;
      11'h9f: data = 24'b111110000011111000000000;
      11'ha0: data = 24'b111111000011111000000000;
      11'ha1: data = 24'b111111000111111000000000;
      11'ha2: data = 24'b111111000111111000000000;
      11'ha3: data = 24'b111111000111111000000000;
      11'ha4: data = 24'b111111000111111000000000;
      11'ha5: data = 24'b111011101110111000000000;
      11'ha6: data = 24'b111011101110111000000000;
      11'ha7: data = 24'b111011101110111000000000;
      11'ha8: data = 24'b111011101110111000000000;
      11'ha9: data = 24'b111011101110111000000000;
      11'haa: data = 24'b111011111100111000000000;
      11'hab: data = 24'b111001111100111000000000;
      11'hac: data = 24'b111001111100111000000000;
      11'had: data = 24'b111001111100111000000000;
      11'hae: data = 24'b111001111000111000000000;
      11'haf: data = 24'b111000111000111000000000;
      11'hb0: data = 24'b000000000000000000000000;
      11'hb1: data = 24'b000000000000000000000000;
      11'hb2: data = 24'b000000000000000000000000;
      11'hb3: data = 24'b000000000000000000000000;
      11'hb4: data = 24'b000000000000000000000000;
      11'hb5: data = 24'b000000000000000000000000;
      11'hb6: data = 24'b000000000000000000000000;
      11'hb7: data = 24'b000000000000000000000000;
      11'hb8: data = 24'b000000000000000000000000;
      11'hb9: data = 24'b000000000000000000000000;
      11'hba: data = 24'b000000000000000000000000;
      11'hbb: data = 24'b000000000000000000000000;
      11'hbc: data = 24'b000000000000000000000000;
      11'hbd: data = 24'b000000000000000000000000;
      11'hbe: data = 24'b000000000000000000000000;
      11'hbf: data = 24'b000000000000000000000000;

      11'hc0: data = 24'b000000000000000000000000;
      11'hc1: data = 24'b000000000000000000000000;
      11'hc2: data = 24'b000000000000000000000000;
      11'hc3: data = 24'b000000000000000000000000;
      11'hc4: data = 24'b000000000000000000000000;
      11'hc5: data = 24'b000000000000000000000000;
      11'hc6: data = 24'b000000000000000000000000;
      11'hc7: data = 24'b000000000000000000000000;
      11'hc8: data = 24'b000000000000000000000000;
      11'hc9: data = 24'b000000000000000000000000;
      11'hca: data = 24'b000000000000000000000000;
      11'hcb: data = 24'b000000000000000000000000;
      11'hcc: data = 24'b000000000000000000000000;
      11'hcd: data = 24'b000000000000000000000000;
      11'hce: data = 24'b000000000000000000000000;
      11'hcf: data = 24'b000000111111000000000000;
      11'hd0: data = 24'b000011111111100000000000;
      11'hd1: data = 24'b000111110011110000000000;
      11'hd2: data = 24'b000111100001110000000000;
      11'hd3: data = 24'b000111100001110000000000;
      11'hd4: data = 24'b001111000001111000000000;
      11'hd5: data = 24'b001111000001111000000000;
      11'hd6: data = 24'b001111111111111000000000;
      11'hd7: data = 24'b001111111111111000000000;
      11'hd8: data = 24'b001111000000000000000000;
      11'hd9: data = 24'b001111000000000000000000;
      11'hda: data = 24'b001111000001111000000000;
      11'hdb: data = 24'b000111100011110000000000;
      11'hdc: data = 24'b000111100011110000000000;
      11'hdd: data = 24'b000111110011110000000000;
      11'hde: data = 24'b000011111111100000000000;
      11'hdf: data = 24'b000001111111000000000000;
      11'he0: data = 24'b000000000000000000000000;
      11'he1: data = 24'b000000000000000000000000;
      11'he2: data = 24'b000000000000000000000000;
      11'he3: data = 24'b000000000000000000000000;
      11'he4: data = 24'b000000000000000000000000;
      11'he5: data = 24'b000000000000000000000000;
      11'he6: data = 24'b000000000000000000000000;
      11'he7: data = 24'b000000000000000000000000;
      11'he8: data = 24'b000000000000000000000000;
      11'he9: data = 24'b000000000000000000000000;
      11'hea: data = 24'b000000000000000000000000;
      11'heb: data = 24'b000000000000000000000000;
      11'hec: data = 24'b000000000000000000000000;
      11'hed: data = 24'b000000000000000000000000;
      11'hee: data = 24'b000000000000000000000000;
      11'hef: data = 24'b000000000000000000000000;

      11'hf0: data = 24'b000000000000000000000000;
      11'hf1: data = 24'b000000000000000000000000;
      11'hf2: data = 24'b000000000000000000000000;
      11'hf3: data = 24'b000000000000000000000000;
      11'hf4: data = 24'b000000000000000000000000;
      11'hf5: data = 24'b000000000000000000000000;
      11'hf6: data = 24'b000000000000000000000000;
      11'hf7: data = 24'b000000000000000000000000;
      11'hf8: data = 24'b000000000000000000000000;
      11'hf9: data = 24'b000000000000000000000000;
      11'hfa: data = 24'b000000000000000000000000;
      11'hfb: data = 24'b000000000000000000000000;
      11'hfc: data = 24'b000000000000000000000000;
      11'hfd: data = 24'b000000000000000000000000;
      11'hfe: data = 24'b000000000000000000000000;
      11'hff: data = 24'b000001111110000000000000;
      11'h100: data = 24'b000111111111100000000000;
      11'h101: data = 24'b000111100111110000000000;
      11'h102: data = 24'b001111000011110000000000;
      11'h103: data = 24'b001111000011110000000000;
      11'h104: data = 24'b001111110000000000000000;
      11'h105: data = 24'b000111111110000000000000;
      11'h106: data = 24'b000011111111100000000000;
      11'h107: data = 24'b000000111111110000000000;
      11'h108: data = 24'b000000000111110000000000;
      11'h109: data = 24'b000000000011111000000000;
      11'h10a: data = 24'b000000000001111000000000;
      11'h10b: data = 24'b001111000001110000000000;
      11'h10c: data = 24'b001111000011110000000000;
      11'h10d: data = 24'b000111100011110000000000;
      11'h10e: data = 24'b000111111111100000000000;
      11'h10f: data = 24'b000001111111000000000000;
      11'h110: data = 24'b000000000000000000000000;
      11'h111: data = 24'b000000000000000000000000;
      11'h112: data = 24'b000000000000000000000000;
      11'h113: data = 24'b000000000000000000000000;
      11'h114: data = 24'b000000000000000000000000;
      11'h115: data = 24'b000000000000000000000000;
      11'h116: data = 24'b000000000000000000000000;
      11'h117: data = 24'b000000000000000000000000;
      11'h118: data = 24'b000000000000000000000000;
      11'h119: data = 24'b000000000000000000000000;
      11'h11a: data = 24'b000000000000000000000000;
      11'h11b: data = 24'b000000000000000000000000;
      11'h11c: data = 24'b000000000000000000000000;
      11'h11d: data = 24'b000000000000000000000000;
      11'h11e: data = 24'b000000000000000000000000;
      11'h11f: data = 24'b000000000000000000000000;

      
      11'h120: data = 24'b000000000000000000000000;
      11'h121: data = 24'b000000000000000000000000;
      11'h122: data = 24'b000000000000000000000000;
      11'h123: data = 24'b000000000000000000000000;
      11'h124: data = 24'b000000000000000000000000;
      11'h125: data = 24'b000000000000000000000000;
      11'h126: data = 24'b000000000000000000000000;
      11'h127: data = 24'b000000000000000000000000;
      11'h128: data = 24'b000000000000000000000000;
      11'h129: data = 24'b000000011100000000000000;
      11'h12a: data = 24'b000000011100000000000000;
      11'h12b: data = 24'b000000111110000000000000;
      11'h12c: data = 24'b000000111110000000000000;
      11'h12d: data = 24'b000001111111000000000000;
      11'h12e: data = 24'b000001111111000000000000;
      11'h12f: data = 24'b000001111111000000000000;
      11'h130: data = 24'b000011110111100000000000;
      11'h131: data = 24'b000011110111100000000000;
      11'h132: data = 24'b000011100111100000000000;
      11'h133: data = 24'b000111100011110000000000;
      11'h134: data = 24'b000111100011110000000000;
      11'h135: data = 24'b000111000001110000000000;
      11'h136: data = 24'b001111000001111000000000;
      11'h137: data = 24'b001111111111111000000000;
      11'h138: data = 24'b001111111111111000000000;
      11'h139: data = 24'b011110000000111100000000;
      11'h13a: data = 24'b011110000000111100000000;
      11'h13b: data = 24'b011110000000111100000000;
      11'h13c: data = 24'b011110000000111100000000;
      11'h13d: data = 24'b011110000000111100000000;
      11'h13e: data = 24'b011110000000111100000000;
      11'h13f: data = 24'b011110000000111100000000;
      11'h140: data = 24'b000000000000000000000000;
      11'h141: data = 24'b000000000000000000000000;
      11'h142: data = 24'b000000000000000000000000;
      11'h143: data = 24'b000000000000000000000000;
      11'h144: data = 24'b000000000000000000000000;
      11'h145: data = 24'b000000000000000000000000;
      11'h146: data = 24'b000000000000000000000000;
      11'h147: data = 24'b000000000000000000000000;
      11'h148: data = 24'b000000000000000000000000;
      11'h149: data = 24'b000000000000000000000000;
      11'h14a: data = 24'b000000000000000000000000;
      11'h14b: data = 24'b000000000000000000000000;
      11'h14c: data = 24'b000000000000000000000000;
      11'h14d: data = 24'b000000000000000000000000;
      11'h14e: data = 24'b000000000000000000000000;
      11'h14f: data = 24'b000000000000000000000000;

      11'h150: data = 24'b000000000000000000000000;
      11'h151: data = 24'b000000000000000000000000;
      11'h152: data = 24'b000000000000000000000000;
      11'h153: data = 24'b000000000000000000000000;
      11'h154: data = 24'b000000000000000000000000;
      11'h155: data = 24'b000000000000000000000000;
      11'h156: data = 24'b000000000000000000000000;
      11'h157: data = 24'b000000000000000000000000;
      11'h158: data = 24'b000000000000000000000000;
      11'h159: data = 24'b000000000000000000000000;
      11'h15a: data = 24'b000011110111100000000000;
      11'h15b: data = 24'b000111111111000000000000;
      11'h15c: data = 24'b001111011111000000000000;
      11'h15d: data = 24'b000000000000000000000000;
      11'h15e: data = 24'b000000000000000000000000;
      11'h15f: data = 24'b011111111110000000000000;
      11'h160: data = 24'b011111111111000000000000;
      11'h161: data = 24'b011111100111100000000000;
      11'h162: data = 24'b011111000111100000000000;
      11'h163: data = 24'b011110000011110000000000;
      11'h164: data = 24'b011110000011110000000000;
      11'h165: data = 24'b011110000011110000000000;
      11'h166: data = 24'b011110000011110000000000;
      11'h167: data = 24'b011110000011110000000000;
      11'h168: data = 24'b011110000011110000000000;
      11'h169: data = 24'b011110000011110000000000;
      11'h16a: data = 24'b011110000011110000000000;
      11'h16b: data = 24'b011110000011110000000000;
      11'h16c: data = 24'b011110000011110000000000;
      11'h16d: data = 24'b011110000011110000000000;
      11'h16e: data = 24'b011110000011110000000000;
      11'h16f: data = 24'b011110000011110000000000;
      11'h170: data = 24'b000000000000000000000000;
      11'h171: data = 24'b000000000000000000000000;
      11'h172: data = 24'b000000000000000000000000;
      11'h173: data = 24'b000000000000000000000000;
      11'h174: data = 24'b000000000000000000000000;
      11'h175: data = 24'b000000000000000000000000;
      11'h176: data = 24'b000000000000000000000000;
      11'h177: data = 24'b000000000000000000000000;
      11'h178: data = 24'b000000000000000000000000;
      11'h179: data = 24'b000000000000000000000000;
      11'h17a: data = 24'b000000000000000000000000;
      11'h17b: data = 24'b000000000000000000000000;
      11'h17c: data = 24'b000000000000000000000000;
      11'h17d: data = 24'b000000000000000000000000;
      11'h17e: data = 24'b000000000000000000000000;
      11'h17f: data = 24'b000000000000000000000000;

      11'h180: data = 24'b000000000000000000000000;
      11'h181: data = 24'b000000000000000000000000;
      11'h182: data = 24'b000000000000000000000000;
      11'h183: data = 24'b000000000000000000000000;
      11'h184: data = 24'b000000000000000000000000;
      11'h185: data = 24'b000000000000000000000000;
      11'h186: data = 24'b000000000000000000000000;
      11'h187: data = 24'b000000000000000000000000;
      11'h188: data = 24'b000000000000000000000000;
      11'h189: data = 24'b000000000000000000000000;
      11'h18a: data = 24'b000000000000000000000000;
      11'h18b: data = 24'b000000000000000000000000;
      11'h18c: data = 24'b000000000000000000000000;
      11'h18d: data = 24'b000000000000000000000000;
      11'h18e: data = 24'b000000000000000000000000;
      11'h18f: data = 24'b000001111111000000000000;
      11'h190: data = 24'b000011111111100000000000;
      11'h191: data = 24'b000111100111110000000000;
      11'h192: data = 24'b001111000001111000000000;
      11'h193: data = 24'b001111000001111000000000;
      11'h194: data = 24'b011110000000111000000000;
      11'h195: data = 24'b011110000000111000000000;
      11'h196: data = 24'b011110000000111000000000;
      11'h197: data = 24'b011110000000111000000000;
      11'h198: data = 24'b011110000000111000000000;
      11'h199: data = 24'b011110000000111000000000;
      11'h19a: data = 24'b011110000001111000000000;
      11'h19b: data = 24'b001111000001111000000000;
      11'h19c: data = 24'b001111000001111000000000;
      11'h19d: data = 24'b000111100111110000000000;
      11'h19e: data = 24'b000011111111100000000000;
      11'h19f: data = 24'b000001111111000000000000;
      11'h1a0: data = 24'b000000000000000000000000;
      11'h1a1: data = 24'b000000000000000000000000;
      11'h1a2: data = 24'b000000000000000000000000;
      11'h1a3: data = 24'b000000000000000000000000;
      11'h1a4: data = 24'b000000000000000000000000;
      11'h1a5: data = 24'b000000000000000000000000;
      11'h1a6: data = 24'b000000000000000000000000;
      11'h1a7: data = 24'b000000000000000000000000;
      11'h1a8: data = 24'b000000000000000000000000;
      11'h1a9: data = 24'b000000000000000000000000;
      11'h1aa: data = 24'b000000000000000000000000;
      11'h1ab: data = 24'b000000000000000000000000;
      11'h1ac: data = 24'b000000000000000000000000;
      11'h1ad: data = 24'b000000000000000000000000;
      11'h1ae: data = 24'b000000000000000000000000;
      11'h1af: data = 24'b000000000000000000000000;

      11'h1b0: data = 24'b000000000000000000000000;
      11'h1b1: data = 24'b000000000000000000000000;
      11'h1b2: data = 24'b000000000000000000000000;
      11'h1b3: data = 24'b000000000000000000000000;
      11'h1b4: data = 24'b000000000000000000000000;
      11'h1b5: data = 24'b000000000000000000000000;
      11'h1b6: data = 24'b000000000000000000000000;
      11'h1b7: data = 24'b000000000000000000000000;
      11'h1b8: data = 24'b000000000000000000000000;
      11'h1b9: data = 24'b000000000000000000000000;
      11'h1ba: data = 24'b000000000000000000000000;
      11'h1bb: data = 24'b000001111110000000000000;
      11'h1bc: data = 24'b000111111111100000000000;
      11'h1bd: data = 24'b001111000111110000000000;
      11'h1be: data = 24'b011110000011110000000000;
      11'h1bf: data = 24'b111100000001111000000000;
      11'h1c0: data = 24'b111100000001111000000000;
      11'h1c1: data = 24'b111000000000110000000000;
      11'h1c2: data = 24'b111000000000000000000000;
      11'h1c3: data = 24'b111000000000000000000000;
      11'h1c4: data = 24'b111000000000000000000000;
      11'h1c5: data = 24'b111000000000000000000000;
      11'h1c6: data = 24'b111000000000000000000000;
      11'h1c7: data = 24'b111000000000000000000000;
      11'h1c8: data = 24'b111000000000111000000000;
      11'h1c9: data = 24'b111000000000111000000000;
      11'h1ca: data = 24'b111100000001111000000000;
      11'h1cb: data = 24'b011100000001111000000000;
      11'h1cc: data = 24'b011110000011110000000000;
      11'h1cd: data = 24'b001111000111110000000000;
      11'h1ce: data = 24'b000111111111100000000000;
      11'h1cf: data = 24'b000011111110000000000000;
      11'h1d0: data = 24'b000000000000000000000000;
      11'h1d1: data = 24'b000000000000000000000000;
      11'h1d2: data = 24'b000000000000000000000000;
      11'h1d3: data = 24'b000000000000000000000000;
      11'h1d4: data = 24'b000000000000000000000000;
      11'h1d5: data = 24'b000000000000000000000000;
      11'h1d6: data = 24'b000000000000000000000000;
      11'h1d7: data = 24'b000000000000000000000000;
      11'h1d8: data = 24'b000000000000000000000000;
      11'h1d9: data = 24'b000000000000000000000000;
      11'h1da: data = 24'b000000000000000000000000;
      11'h1db: data = 24'b000000000000000000000000;
      11'h1dc: data = 24'b000000000000000000000000;
      11'h1dd: data = 24'b000000000000000000000000;
      11'h1de: data = 24'b000000000000000000000000;
      11'h1df: data = 24'b000000000000000000000000;

      11'h1e0: data = 24'b000000000000000000000000;
      11'h1e1: data = 24'b000000000000000000000000;
      11'h1e2: data = 24'b000000000000000000000000;
      11'h1e3: data = 24'b000000000000000000000000;
      11'h1e4: data = 24'b000000000000000000000000;
      11'h1e5: data = 24'b000000000000000000000000;
      11'h1e6: data = 24'b000000000000000000000000;
      11'h1e7: data = 24'b000000000000000000000000;
      11'h1e8: data = 24'b000000000000000000000000;
      11'h1e9: data = 24'b000000000000000000000000;
      11'h1ea: data = 24'b000000000000000000000000;
      11'h1eb: data = 24'b000000000000000000000000;
      11'h1ec: data = 24'b000000000000000000000000;
      11'h1ed: data = 24'b000000000000000000000000;
      11'h1ee: data = 24'b000000000000000000000000;
      11'h1ef: data = 24'b000001101110000000000000;
      11'h1f0: data = 24'b000001111111000000000000;
      11'h1f1: data = 24'b000001111111000000000000;
      11'h1f2: data = 24'b000001111011000000000000;
      11'h1f3: data = 24'b000001111011000000000000;
      11'h1f4: data = 24'b000001111011000000000000;
      11'h1f5: data = 24'b000001110000000000000000;
      11'h1f6: data = 24'b000001110000000000000000;
      11'h1f7: data = 24'b000001110000000000000000;
      11'h1f8: data = 24'b000001110000000000000000;
      11'h1f9: data = 24'b000001110000000000000000;
      11'h1fa: data = 24'b000001110000000000000000;
      11'h1fb: data = 24'b000001110000000000000000;
      11'h1fc: data = 24'b000001110000000000000000;
      11'h1fd: data = 24'b000001110000000000000000;
      11'h1fe: data = 24'b000001110000000000000000;
      11'h1ff: data = 24'b000001110000000000000000;
      11'h200: data = 24'b000000000000000000000000;
      11'h201: data = 24'b000000000000000000000000;
      11'h202: data = 24'b000000000000000000000000;
      11'h203: data = 24'b000000000000000000000000;
      11'h204: data = 24'b000000000000000000000000;
      11'h205: data = 24'b000000000000000000000000;
      11'h206: data = 24'b000000000000000000000000;
      11'h207: data = 24'b000000000000000000000000;
      11'h208: data = 24'b000000000000000000000000;
      11'h209: data = 24'b000000000000000000000000;
      11'h20a: data = 24'b000000000000000000000000;
      11'h20b: data = 24'b000000000000000000000000;
      11'h20c: data = 24'b000000000000000000000000;
      11'h20d: data = 24'b000000000000000000000000;
      11'h20e: data = 24'b000000000000000000000000;
      11'h20f: data = 24'b000000000000000000000000;

      11'h210: data = 24'b000000000000000000000000;
      11'h211: data = 24'b000000000000000000000000;
      11'h212: data = 24'b000000000000000000000000;
      11'h213: data = 24'b000000000000000000000000;
      11'h214: data = 24'b000000000000000000000000;
      11'h215: data = 24'b000000000000000000000000;
      11'h216: data = 24'b000000000000000000000000;
      11'h217: data = 24'b000000000000000000000000;
      11'h218: data = 24'b000000000000000000000000;
      11'h219: data = 24'b000000000000000000000000;
      11'h21a: data = 24'b000000000000000000000000;
      11'h21b: data = 24'b000000000000000000000000;
      11'h21c: data = 24'b000000000000000000000000;
      11'h21d: data = 24'b000000000000000000000000;
      11'h21e: data = 24'b000000000000000000000000;
      11'h21f: data = 24'b011110111111000000000000;
      11'h220: data = 24'b011111111111110000000000;
      11'h221: data = 24'b011111111111111000000000;
      11'h222: data = 24'b011111110011111000000000;
      11'h223: data = 24'b011111000001111000000000;
      11'h224: data = 24'b011111000001111000000000;
      11'h225: data = 24'b011111000001111000000000;
      11'h226: data = 24'b011111000001111000000000;
      11'h227: data = 24'b011110000001111000000000;
      11'h228: data = 24'b011110000001111000000000;
      11'h229: data = 24'b011110000001111000000000;
      11'h22a: data = 24'b011110000001111000000000;
      11'h22b: data = 24'b011110000001111000000000;
      11'h22c: data = 24'b011110000001111000000000;
      11'h22d: data = 24'b011110000001111000000000;
      11'h22e: data = 24'b011110000001111000000000;
      11'h22f: data = 24'b011110000001111000000000;
      11'h230: data = 24'b000000000000000000000000;
      11'h231: data = 24'b000000000000000000000000;
      11'h232: data = 24'b000000000000000000000000;
      11'h233: data = 24'b000000000000000000000000;
      11'h234: data = 24'b000000000000000000000000;
      11'h235: data = 24'b000000000000000000000000;
      11'h236: data = 24'b000000000000000000000000;
      11'h237: data = 24'b000000000000000000000000;
      11'h238: data = 24'b000000000000000000000000;
      11'h239: data = 24'b000000000000000000000000;
      11'h23a: data = 24'b000000000000000000000000;
      11'h23b: data = 24'b000000000000000000000000;
      11'h23c: data = 24'b000000000000000000000000;
      11'h23d: data = 24'b000000000000000000000000;
      11'h23e: data = 24'b000000000000000000000000;
      11'h23f: data = 24'b000000000000000000000000;

      11'h240: data = 24'b000000000000000000000000;
      11'h241: data = 24'b000000000000000000000000;
      11'h242: data = 24'b000000000000000000000000;
      11'h243: data = 24'b000000000000000000000000;
      11'h244: data = 24'b000000000000000000000000;
      11'h245: data = 24'b000000000000000000000000;
      11'h246: data = 24'b000000000000000000000000;
      11'h247: data = 24'b000000000000000000000000;
      11'h248: data = 24'b000000000000000000000000;
      11'h249: data = 24'b000000000000000000000000;
      11'h24a: data = 24'b000000000000000000000000;
      11'h24b: data = 24'b000000000000000000000000;
      11'h24c: data = 24'b000000000000000000000000;
      11'h24d: data = 24'b000000000000000000000000;
      11'h24e: data = 24'b000000000000000000000000;
      11'h24f: data = 24'b111111110011111000000000;
      11'h250: data = 24'b111111111111111100000000;
      11'h251: data = 24'b111100111110111100000000;
      11'h252: data = 24'b111100111100011100000000;
      11'h253: data = 24'b111100111100011100000000;
      11'h254: data = 24'b111000111100011100000000;
      11'h255: data = 24'b111000111100011100000000;
      11'h256: data = 24'b111000111100011100000000;
      11'h257: data = 24'b111000111100011100000000;
      11'h258: data = 24'b111000111100011100000000;
      11'h259: data = 24'b111000111100011100000000;
      11'h25a: data = 24'b111000111100011100000000;
      11'h25b: data = 24'b111000111100011100000000;
      11'h25c: data = 24'b111000111100011100000000;
      11'h25d: data = 24'b111000111100011100000000;
      11'h25e: data = 24'b111000111100011100000000;
      11'h25f: data = 24'b111000111100011100000000;
      11'h260: data = 24'b000000000000000000000000;
      11'h261: data = 24'b000000000000000000000000;
      11'h262: data = 24'b000000000000000000000000;
      11'h263: data = 24'b000000000000000000000000;
      11'h264: data = 24'b000000000000000000000000;
      11'h265: data = 24'b000000000000000000000000;
      11'h266: data = 24'b000000000000000000000000;
      11'h267: data = 24'b000000000000000000000000;
      11'h268: data = 24'b000000000000000000000000;
      11'h269: data = 24'b000000000000000000000000;
      11'h26a: data = 24'b000000000000000000000000;
      11'h26b: data = 24'b000000000000000000000000;
      11'h26c: data = 24'b000000000000000000000000;
      11'h26d: data = 24'b000000000000000000000000;
      11'h26e: data = 24'b000000000000000000000000;
      11'h26f: data = 24'b000000000000000000000000;

      11'h270: data = 24'b000000000000000000000000;
      11'h271: data = 24'b000000000000000000000000;
      11'h272: data = 24'b000000000000000000000000;
      11'h273: data = 24'b000000000000000000000000;
      11'h274: data = 24'b000000000000000000000000;
      11'h275: data = 24'b000000000000000000000000;
      11'h276: data = 24'b000000000000000000000000;
      11'h277: data = 24'b000000000000000000000000;
      11'h278: data = 24'b000000000000000000000000;
      11'h279: data = 24'b000000000000000000000000;
      11'h27a: data = 24'b000000011000000000000000;
      11'h27b: data = 24'b000000111000000000000000;
      11'h27c: data = 24'b000001111000000000000000;
      11'h27d: data = 24'b000001111000000000000000;
      11'h27e: data = 24'b000001111000000000000000;
      11'h27f: data = 24'b000011111110000000000000;
      11'h280: data = 24'b000011111110000000000000;
      11'h281: data = 24'b000001111000000000000000;
      11'h282: data = 24'b000001111000000000000000;
      11'h283: data = 24'b000001111000000000000000;
      11'h284: data = 24'b000001111000000000000000;
      11'h285: data = 24'b000001111000000000000000;
      11'h286: data = 24'b000001111000000000000000;
      11'h287: data = 24'b000001111000000000000000;
      11'h288: data = 24'b000001111000000000000000;
      11'h289: data = 24'b000001111000000000000000;
      11'h28a: data = 24'b000001111000000000000000;
      11'h28b: data = 24'b000001111000000000000000;
      11'h28c: data = 24'b000001111000000000000000;
      11'h28d: data = 24'b000001111000000000000000;
      11'h28e: data = 24'b000000111111000000000000;
      11'h28f: data = 24'b000000011111000000000000;
      11'h290: data = 24'b000000000000000000000000;
      11'h291: data = 24'b000000000000000000000000;
      11'h292: data = 24'b000000000000000000000000;
      11'h293: data = 24'b000000000000000000000000;
      11'h294: data = 24'b000000000000000000000000;
      11'h295: data = 24'b000000000000000000000000;
      11'h296: data = 24'b000000000000000000000000;
      11'h297: data = 24'b000000000000000000000000;
      11'h298: data = 24'b000000000000000000000000;
      11'h299: data = 24'b000000000000000000000000;
      11'h29a: data = 24'b000000000000000000000000;
      11'h29b: data = 24'b000000000000000000000000;
      11'h29c: data = 24'b000000000000000000000000;
      11'h29d: data = 24'b000000000000000000000000;
      11'h29e: data = 24'b000000000000000000000000;
      11'h29f: data = 24'b000000000000000000000000;

      11'h2a0: data = 24'b000000000000000000000000;
      11'h2a1: data = 24'b000000000000000000000000;
      11'h2a2: data = 24'b000000000000000000000000;
      11'h2a3: data = 24'b000000000000000000000000;
      11'h2a4: data = 24'b000000000000000000000000;
      11'h2a5: data = 24'b000000000000000000000000;
      11'h2a6: data = 24'b000000000000000000000000;
      11'h2a7: data = 24'b000000000000000000000000;
      11'h2a8: data = 24'b000000000000000000000000;
      11'h2a9: data = 24'b111111111111000000000000;
      11'h2aa: data = 24'b111111111111110000000000;
      11'h2ab: data = 24'b111100000011110000000000;
      11'h2ac: data = 24'b111100000001111000000000;
      11'h2ad: data = 24'b111100000001111000000000;
      11'h2ae: data = 24'b111100000001111000000000;
      11'h2af: data = 24'b111100000001111000000000;
      11'h2b0: data = 24'b111100000001111000000000;
      11'h2b1: data = 24'b111100000001111000000000;
      11'h2b2: data = 24'b111100000011110000000000;
      11'h2b3: data = 24'b111111111111100000000000;
      11'h2b4: data = 24'b111111111100000000000000;
      11'h2b5: data = 24'b111100011110000000000000;
      11'h2b6: data = 24'b111100001111000000000000;
      11'h2b7: data = 24'b111100000111100000000000;
      11'h2b8: data = 24'b111100000111100000000000;
      11'h2b9: data = 24'b111100000011110000000000;
      11'h2ba: data = 24'b111100000011110000000000;
      11'h2bb: data = 24'b111100000011110000000000;
      11'h2bc: data = 24'b111100000001111000000000;
      11'h2bd: data = 24'b111100000001111000000000;
      11'h2be: data = 24'b111100000000111000000000;
      11'h2bf: data = 24'b111100000000111000000000;
      11'h2c0: data = 24'b000000000000000000000000;
      11'h2c1: data = 24'b000000000000000000000000;
      11'h2c2: data = 24'b000000000000000000000000;
      11'h2c3: data = 24'b000000000000000000000000;
      11'h2c4: data = 24'b000000000000000000000000;
      11'h2c5: data = 24'b000000000000000000000000;
      11'h2c6: data = 24'b000000000000000000000000;
      11'h2c7: data = 24'b000000000000000000000000;
      11'h2c8: data = 24'b000000000000000000000000;
      11'h2c9: data = 24'b000000000000000000000000;
      11'h2ca: data = 24'b000000000000000000000000;
      11'h2cb: data = 24'b000000000000000000000000;
      11'h2cc: data = 24'b000000000000000000000000;
      11'h2cd: data = 24'b000000000000000000000000;
      11'h2ce: data = 24'b000000000000000000000000;
      11'h2cf: data = 24'b000000000000000000000000;

      11'h2d0: data = 24'b000000000000000000000000;
      11'h2d1: data = 24'b000000000000000000000000;
      11'h2d2: data = 24'b000000000000000000000000;
      11'h2d3: data = 24'b000000000000000000000000;
      11'h2d4: data = 24'b000000000000000000000000;
      11'h2d5: data = 24'b000000000000000000000000;
      11'h2d6: data = 24'b000000000000000000000000;
      11'h2d7: data = 24'b000000000000000000000000;
      11'h2d8: data = 24'b000000000000000000000000;
      11'h2d9: data = 24'b000000000000000000000000;
      11'h2da: data = 24'b000000000000000000000000;
      11'h2db: data = 24'b000000000000000000000000;
      11'h2dc: data = 24'b000000000000000000000000;
      11'h2dd: data = 24'b000000000000000000000000;
      11'h2de: data = 24'b000000000000000000000000;
      11'h2df: data = 24'b000011111101110000000000;
      11'h2e0: data = 24'b000111111111110000000000;
      11'h2e1: data = 24'b001111000111110000000000;
      11'h2e2: data = 24'b011110000111110000000000;
      11'h2e3: data = 24'b011110000011110000000000;
      11'h2e4: data = 24'b011110000011110000000000;
      11'h2e5: data = 24'b011110000011110000000000;
      11'h2e6: data = 24'b011110000011110000000000;
      11'h2e7: data = 24'b011110000111110000000000;
      11'h2e8: data = 24'b001111000111110000000000;
      11'h2e9: data = 24'b001111001111110000000000;
      11'h2ea: data = 24'b000111111111110000000000;
      11'h2eb: data = 24'b000000000011110000000000;
      11'h2ec: data = 24'b011110000011100000000000;
      11'h2ed: data = 24'b011110000111100000000000;
      11'h2ee: data = 24'b001111111111100000000000;
      11'h2ef: data = 24'b000011111111000000000000;
      11'h2f0: data = 24'b000000000000000000000000;
      11'h2f1: data = 24'b000000000000000000000000;
      11'h2f2: data = 24'b000000000000000000000000;
      11'h2f3: data = 24'b000000000000000000000000;
      11'h2f4: data = 24'b000000000000000000000000;
      11'h2f5: data = 24'b000000000000000000000000;
      11'h2f6: data = 24'b000000000000000000000000;
      11'h2f7: data = 24'b000000000000000000000000;
      11'h2f8: data = 24'b000000000000000000000000;
      11'h2f9: data = 24'b000000000000000000000000;
      11'h2fa: data = 24'b000000000000000000000000;
      11'h2fb: data = 24'b000000000000000000000000;
      11'h2fc: data = 24'b000000000000000000000000;
      11'h2fd: data = 24'b000000000000000000000000;
      11'h2fe: data = 24'b000000000000000000000000;
      11'h2ff: data = 24'b000000000000000000000000;

      11'h300: data = 24'b000000000000000000000000;
      11'h301: data = 24'b000000000000000000000000;
      11'h302: data = 24'b000000000000000000000000;
      11'h303: data = 24'b000000000000000000000000;
      11'h304: data = 24'b000000000000000000000000;
      11'h305: data = 24'b000000000000000000000000;
      11'h306: data = 24'b000000000000000000000000;
      11'h307: data = 24'b000000000000000000000000;
      11'h308: data = 24'b000000000000000000000000;
      11'h309: data = 24'b000000000000000000000000;
      11'h30a: data = 24'b000000000000000000000000;
      11'h30b: data = 24'b111100000001111000000000;
      11'h30c: data = 24'b111100000001111000000000;
      11'h30d: data = 24'b111100000001111000000000;
      11'h30e: data = 24'b111100000001111000000000;
      11'h30f: data = 24'b111100000001111000000000;
      11'h310: data = 24'b111100000001111000000000;
      11'h311: data = 24'b111100000001111000000000;
      11'h312: data = 24'b111100000001111000000000;
      11'h313: data = 24'b111100000001111000000000;
      11'h314: data = 24'b111111111111111000000000;
      11'h315: data = 24'b111111111111111000000000;
      11'h316: data = 24'b111100000001111000000000;
      11'h317: data = 24'b111100000001111000000000;
      11'h318: data = 24'b111100000001111000000000;
      11'h319: data = 24'b111100000001111000000000;
      11'h31a: data = 24'b111100000001111000000000;
      11'h31b: data = 24'b111100000001111000000000;
      11'h31c: data = 24'b111100000001111000000000;
      11'h31d: data = 24'b111100000001111000000000;
      11'h31e: data = 24'b111100000001111000000000;
      11'h31f: data = 24'b111100000001111000000000;
      11'h320: data = 24'b000000000000000000000000;
      11'h321: data = 24'b000000000000000000000000;
      11'h322: data = 24'b000000000000000000000000;
      11'h323: data = 24'b000000000000000000000000;
      11'h324: data = 24'b000000000000000000000000;
      11'h325: data = 24'b000000000000000000000000;
      11'h326: data = 24'b000000000000000000000000;
      11'h327: data = 24'b000000000000000000000000;
      11'h328: data = 24'b000000000000000000000000;
      11'h329: data = 24'b000000000000000000000000;
      11'h32a: data = 24'b000000000000000000000000;
      11'h32b: data = 24'b000000000000000000000000;
      11'h32c: data = 24'b000000000000000000000000;
      11'h32d: data = 24'b000000000000000000000000;
      11'h32e: data = 24'b000000000000000000000000;
      11'h32f: data = 24'b000000000000000000000000;

      11'h330: data = 24'b000000000000000000000000;
      11'h331: data = 24'b000000000000000000000000;
      11'h332: data = 24'b000000000000000000000000;
      11'h333: data = 24'b000000000000000000000000;
      11'h334: data = 24'b000000000000000000000000;
      11'h335: data = 24'b000000000000000000000000;
      11'h336: data = 24'b000000000000000000000000;
      11'h337: data = 24'b000000000000000000000000;
      11'h338: data = 24'b000000000000000000000000;
      11'h339: data = 24'b000000000000000000000000;
      11'h33a: data = 24'b000000000000000000000000;
      11'h33b: data = 24'b000011111111000000000000;
      11'h33c: data = 24'b000111111111100000000000;
      11'h33d: data = 24'b001111000011110000000000;
      11'h33e: data = 24'b011110000001111000000000;
      11'h33f: data = 24'b011110000001111000000000;
      11'h340: data = 24'b011110000000000000000000;
      11'h341: data = 24'b011110000000000000000000;
      11'h342: data = 24'b011111000000000000000000;
      11'h343: data = 24'b001111110000000000000000;
      11'h344: data = 24'b000111111110000000000000;
      11'h345: data = 24'b000011111111100000000000;
      11'h346: data = 24'b000000011111110000000000;
      11'h347: data = 24'b000000000011111000000000;
      11'h348: data = 24'b000000000001111000000000;
      11'h349: data = 24'b000000000000111000000000;
      11'h34a: data = 24'b111100000000111000000000;
      11'h34b: data = 24'b011100000000111000000000;
      11'h34c: data = 24'b011110000001111000000000;
      11'h34d: data = 24'b011111000011110000000000;
      11'h34e: data = 24'b001111111111100000000000;
      11'h34f: data = 24'b000011111111000000000000;
      11'h350: data = 24'b000000000000000000000000;
      11'h351: data = 24'b000000000000000000000000;
      11'h352: data = 24'b000000000000000000000000;
      11'h353: data = 24'b000000000000000000000000;
      11'h354: data = 24'b000000000000000000000000;
      11'h355: data = 24'b000000000000000000000000;
      11'h356: data = 24'b000000000000000000000000;
      11'h357: data = 24'b000000000000000000000000;
      11'h358: data = 24'b000000000000000000000000;
      11'h359: data = 24'b000000000000000000000000;
      11'h35a: data = 24'b000000000000000000000000;
      11'h35b: data = 24'b000000000000000000000000;
      11'h35c: data = 24'b000000000000000000000000;
      11'h35d: data = 24'b000000000000000000000000;
      11'h35e: data = 24'b000000000000000000000000;
      11'h35f: data = 24'b000000000000000000000000;

      11'h360: data = 24'b000000000000000000000000;
      11'h361: data = 24'b000000000000000000000000;
      11'h362: data = 24'b000000000000000000000000;
      11'h363: data = 24'b000000000000000000000000;
      11'h364: data = 24'b000000000000000000000000;
      11'h365: data = 24'b000000000000000000000000;
      11'h366: data = 24'b000000000000000000000000;
      11'h367: data = 24'b000000000000000000000000;
      11'h368: data = 24'b000000000000000000000000;
      11'h369: data = 24'b000000000000000000000000;
      11'h36a: data = 24'b000000000000000000000000;
      11'h36b: data = 24'b000000000000000000000000;
      11'h36c: data = 24'b000000000000000000000000;
      11'h36d: data = 24'b000000000000000000000000;
      11'h36e: data = 24'b000000000000000000000000;
      11'h36f: data = 24'b000000000000000000000000;
      11'h370: data = 24'b011111000000000000011110;
      11'h371: data = 24'b011111000000000000011110;
      11'h372: data = 24'b011111000000000000011110;
      11'h373: data = 24'b011111000000000000011110;
      11'h374: data = 24'b011111000000000000011110;
      11'h375: data = 24'b011111000000000000011110;
      11'h376: data = 24'b011111000000000000011110;
      11'h377: data = 24'b011111000000000000011110;
      11'h378: data = 24'b011111000000000000011110;
      11'h379: data = 24'b011111000000000000011110;
      11'h37a: data = 24'b011111000000000000011110;
      11'h37b: data = 24'b011111000000000000011110;
      11'h37c: data = 24'b011111000000000000011110;
      11'h37d: data = 24'b011111000000000000011110;
      11'h37e: data = 24'b011111111111111111111110;
      11'h37f: data = 24'b011111111111111111111110;
      11'h380: data = 24'b011111111111111111111110;
      11'h381: data = 24'b011111000000000000011110;
      11'h382: data = 24'b011111000000000000011110;
      11'h383: data = 24'b011111000000000000011110;
      11'h384: data = 24'b011111000000000000011110;
      11'h385: data = 24'b011111000000000000011110;
      11'h386: data = 24'b011111000000000000011110;
      11'h387: data = 24'b011111000000000000011110;
      11'h388: data = 24'b011111000000000000011110;
      11'h389: data = 24'b011111000000000000011110;
      11'h38a: data = 24'b011111000000000000011110;
      11'h38b: data = 24'b011111000000000000011110;
      11'h38c: data = 24'b011111000000000000011110;
      11'h38d: data = 24'b011111000000000000011110;
      11'h38e: data = 24'b011111000000000000011110;
      11'h38f: data = 24'b011111000000000000011110;

      11'h390: data = 24'b000000000000000000000000;
      11'h391: data = 24'b000000000000000000000000;
      11'h392: data = 24'b000000000000000000000000;
      11'h393: data = 24'b000000000000000000000000;
      11'h394: data = 24'b000000000000000000000000;
      11'h395: data = 24'b000000000000000000000000;
      11'h396: data = 24'b000000000000000000000000;
      11'h397: data = 24'b000000000000000000000000;
      11'h398: data = 24'b000000000000000000000000;
      11'h399: data = 24'b000000000000000000000000;
      11'h39a: data = 24'b000000000000000000000000;
      11'h39b: data = 24'b000000000000000000000000;
      11'h39c: data = 24'b000000000000000000000000;
      11'h39d: data = 24'b000000000000000000000000;
      11'h39e: data = 24'b000000000000000000000000;
      11'h39f: data = 24'b000000000000000000000000;
      11'h3a0: data = 24'b000000000000000000000000;
      11'h3a1: data = 24'b000000000000000000000000;
      11'h3a2: data = 24'b000000000000000000000000;
      11'h3a3: data = 24'b000000000000000000000000;
      11'h3a4: data = 24'b000000011111111000000000;
      11'h3a5: data = 24'b000001111111111110000000;
      11'h3a6: data = 24'b000011111111111111000000;
      11'h3a7: data = 24'b000111111111111111100000;
      11'h3a8: data = 24'b000111111100011111110000;
      11'h3a9: data = 24'b001111110000001111110000;
      11'h3aa: data = 24'b001111100000000111111000;
      11'h3ab: data = 24'b011111100000000011111000;
      11'h3ac: data = 24'b011111000000000011111100;
      11'h3ad: data = 24'b011111000000000011111100;
      11'h3ae: data = 24'b011111000000000001111100;
      11'h3af: data = 24'b011111000000000001111100;
      11'h3b0: data = 24'b011111000000000001111100;
      11'h3b1: data = 24'b111111000000000001111100;
      11'h3b2: data = 24'b111111000000000001111100;
      11'h3b3: data = 24'b011111000000000001111100;
      11'h3b4: data = 24'b011111000000000001111100;
      11'h3b5: data = 24'b011111000000000001111100;
      11'h3b6: data = 24'b011111000000000011111100;
      11'h3b7: data = 24'b011111000000000011111100;
      11'h3b8: data = 24'b011111100000000011111000;
      11'h3b9: data = 24'b001111100000000111111000;
      11'h3ba: data = 24'b001111110000001111110000;
      11'h3bb: data = 24'b000111111100011111110000;
      11'h3bc: data = 24'b000111111111111111100000;
      11'h3bd: data = 24'b000011111111111111000000;
      11'h3be: data = 24'b000000111111111110000000;
      11'h3bf: data = 24'b000000001111111000000000;

      11'h3c0: data = 24'b000000000000000000000000;
      11'h3c1: data = 24'b000000000000000000000000;
      11'h3c2: data = 24'b000000000000000000000000;
      11'h3c3: data = 24'b000000000000000000000000;
      11'h3c4: data = 24'b000000000000000000000000;
      11'h3c5: data = 24'b000000000000000000000000;
      11'h3c6: data = 24'b000000000000000000000000;
      11'h3c7: data = 24'b000000000000000000000000;
      11'h3c8: data = 24'b000000000000000000000000;
      11'h3c9: data = 24'b000000000000000000000000;
      11'h3ca: data = 24'b000000000000000000000000;
      11'h3cb: data = 24'b000000000000000000000000;
      11'h3cc: data = 24'b000000000000000000000000;
      11'h3cd: data = 24'b000000000000000000000000;
      11'h3ce: data = 24'b000000000000000000000000;
      11'h3cf: data = 24'b000000000000000000000000;
      11'h3d0: data = 24'b000000000000000000000000;
      11'h3d1: data = 24'b000000000000000000000000;
      11'h3d2: data = 24'b000000000000000000000000;
      11'h3d3: data = 24'b000000000000000000000000;
      11'h3d4: data = 24'b000000000000000000000000;
      11'h3d5: data = 24'b000000000000001111110000;
      11'h3d6: data = 24'b000000001111111111111000;
      11'h3d7: data = 24'b000000001111111111111000;
      11'h3d8: data = 24'b000000001111111111111000;
      11'h3d9: data = 24'b000000001111111100110000;
      11'h3da: data = 24'b000000001111111000000000;
      11'h3db: data = 24'b000000001111110000000000;
      11'h3dc: data = 24'b000000001111110000000000;
      11'h3dd: data = 24'b000000001111110000000000;
      11'h3de: data = 24'b000000001111100000000000;
      11'h3df: data = 24'b000000001111100000000000;
      11'h3e0: data = 24'b000000001111100000000000;
      11'h3e1: data = 24'b000000001111100000000000;
      11'h3e2: data = 24'b000000001111100000000000;
      11'h3e3: data = 24'b000000001111100000000000;
      11'h3e4: data = 24'b000000001111100000000000;
      11'h3e5: data = 24'b000000001111100000000000;
      11'h3e6: data = 24'b000000001111100000000000;
      11'h3e7: data = 24'b000000001111100000000000;
      11'h3e8: data = 24'b000000001111100000000000;
      11'h3e9: data = 24'b000000001111100000000000;
      11'h3ea: data = 24'b000000001111100000000000;
      11'h3eb: data = 24'b000000001111100000000000;
      11'h3ec: data = 24'b000000001111100000000000;
      11'h3ed: data = 24'b000000001111100000000000;
      11'h3ee: data = 24'b000000001111100000000000;
      11'h3ef: data = 24'b000000001111100000000000;

      11'h3f0: data = 24'b000000000000000000000000;
      11'h3f1: data = 24'b000000000000000000000000;
      11'h3f2: data = 24'b000000000000000000000000;
      11'h3f3: data = 24'b000000000000000000000000;
      11'h3f4: data = 24'b000000000000000000000000;
      11'h3f5: data = 24'b000000000000000000000000;
      11'h3f6: data = 24'b000000000000000000000000;
      11'h3f7: data = 24'b000000000000000000000000;
      11'h3f8: data = 24'b000000000000000000000000;
      11'h3f9: data = 24'b000000000000000000000000;
      11'h3fa: data = 24'b000000000000000000000000;
      11'h3fb: data = 24'b000000000000000000000000;
      11'h3fc: data = 24'b000000000000000000000000;
      11'h3fd: data = 24'b000000000000000000000000;
      11'h3fe: data = 24'b000000000000000000000000;
      11'h3ff: data = 24'b000000000000000000000000;
      11'h400: data = 24'b000000000000000000000000;
      11'h401: data = 24'b000000000000000000000000;
      11'h402: data = 24'b000000000000000000000000;
      11'h403: data = 24'b000000000000000000000000;
      11'h404: data = 24'b000000000000000000000000;
      11'h405: data = 24'b000000011111111100000000;
      11'h406: data = 24'b000001111111111111000000;
      11'h407: data = 24'b000111111111111111100000;
      11'h408: data = 24'b000111111111111111110000;
      11'h409: data = 24'b001111111000011111110000;
      11'h40a: data = 24'b001111110000000111110000;
      11'h40b: data = 24'b011111100000000111111000;
      11'h40c: data = 24'b000111100000000011111000;
      11'h40d: data = 24'b000000000000000011111000;
      11'h40e: data = 24'b000000000000000011111000;
      11'h40f: data = 24'b000000000000000111111000;
      11'h410: data = 24'b000000000001111111111000;
      11'h411: data = 24'b000000011111111111111000;
      11'h412: data = 24'b000011111111111111111000;
      11'h413: data = 24'b000111111111111111111000;
      11'h414: data = 24'b001111111111100011111000;
      11'h415: data = 24'b011111111000000011111000;
      11'h416: data = 24'b011111100000000011111000;
      11'h417: data = 24'b011111000000000111111000;
      11'h418: data = 24'b011111000000000111111000;
      11'h419: data = 24'b011111000000000111111000;
      11'h41a: data = 24'b011111000000001111111000;
      11'h41b: data = 24'b011111100000011111111000;
      11'h41c: data = 24'b011111110000111111111000;
      11'h41d: data = 24'b001111111111111111111000;
      11'h41e: data = 24'b001111111111111111111000;
      11'h41f: data = 24'b000111111111110001111100;

      11'h420: data = 24'b000000000000000000000000;
      11'h421: data = 24'b000000000000000000000000;
      11'h422: data = 24'b000000000000000000000000;
      11'h423: data = 24'b000000000000000000000000;
      11'h424: data = 24'b000000000000000000000000;
      11'h425: data = 24'b000000000000000000000000;
      11'h426: data = 24'b000000000000000000000000;
      11'h427: data = 24'b000000000000000000000000;
      11'h428: data = 24'b000000000000000000000000;
      11'h429: data = 24'b000000001111111000000000;
      11'h42a: data = 24'b000000111111111110000000;
      11'h42b: data = 24'b000001111111111111000000;
      11'h42c: data = 24'b000011111111111111000000;
      11'h42d: data = 24'b000011111100111111100000;
      11'h42e: data = 24'b000111111000001111110000;
      11'h42f: data = 24'b000111110000000111110000;
      11'h430: data = 24'b001111110000000111110000;
      11'h431: data = 24'b001111100000000111111000;
      11'h432: data = 24'b001111100000000011111000;
      11'h433: data = 24'b001111100000000011111000;
      11'h434: data = 24'b011111100000000011111000;
      11'h435: data = 24'b011111000000000011111000;
      11'h436: data = 24'b011111000000000011111100;
      11'h437: data = 24'b011111000000000011111100;
      11'h438: data = 24'b011111000000000011111100;
      11'h439: data = 24'b011111000000000001111100;
      11'h43a: data = 24'b011111000000000001111100;
      11'h43b: data = 24'b011111000000000001111100;
      11'h43c: data = 24'b011111000000000001111100;
      11'h43d: data = 24'b011111000000000001111100;
      11'h43e: data = 24'b011111000000000001111100;
      11'h43f: data = 24'b011111000000000001111100;
      11'h440: data = 24'b011111000000000011111100;
      11'h441: data = 24'b011111000000000011111100;
      11'h442: data = 24'b011111000000000011111000;
      11'h443: data = 24'b011111000000000011111000;
      11'h444: data = 24'b011111100000000011111000;
      11'h445: data = 24'b001111100000000011111000;
      11'h446: data = 24'b001111100000000011111000;
      11'h447: data = 24'b001111100000000111111000;
      11'h448: data = 24'b001111110000000111110000;
      11'h449: data = 24'b000111110000000111110000;
      11'h44a: data = 24'b000111111000001111110000;
      11'h44b: data = 24'b000011111100011111100000;
      11'h44c: data = 24'b000011111111111111000000;
      11'h44d: data = 24'b000001111111111111000000;
      11'h44e: data = 24'b000000111111111110000000;
      11'h44f: data = 24'b000000001111111000000000;

      11'h450: data = 24'b000000000000000000000000;
      11'h451: data = 24'b000000000000000000000000;
      11'h452: data = 24'b000000000000000000000000;
      11'h453: data = 24'b000000000000000000000000;
      11'h454: data = 24'b000000000000000000000000;
      11'h455: data = 24'b000000000000000000000000;
      11'h456: data = 24'b000000000000000000000000;
      11'h457: data = 24'b000000000000000000000000;
      11'h458: data = 24'b000000000000000000000000;
      11'h459: data = 24'b000000000000000000000000;
      11'h45a: data = 24'b000000000000000000000000;
      11'h45b: data = 24'b000000000000111100000000;
      11'h45c: data = 24'b000000000000111100000000;
      11'h45d: data = 24'b000000000001111100000000;
      11'h45e: data = 24'b000000000011111100000000;
      11'h45f: data = 24'b000000000011111100000000;
      11'h460: data = 24'b000000000111111100000000;
      11'h461: data = 24'b000000001111111100000000;
      11'h462: data = 24'b000000011111111100000000;
      11'h463: data = 24'b000000111111111100000000;
      11'h464: data = 24'b000011111111111100000000;
      11'h465: data = 24'b000011111101111100000000;
      11'h466: data = 24'b000011111001111100000000;
      11'h467: data = 24'b000011100001111100000000;
      11'h468: data = 24'b000011000001111100000000;
      11'h469: data = 24'b000000000001111100000000;
      11'h46a: data = 24'b000000000001111100000000;
      11'h46b: data = 24'b000000000001111100000000;
      11'h46c: data = 24'b000000000001111100000000;
      11'h46d: data = 24'b000000000001111100000000;
      11'h46e: data = 24'b000000000001111100000000;
      11'h46f: data = 24'b000000000001111100000000;
      11'h470: data = 24'b000000000001111100000000;
      11'h471: data = 24'b000000000001111100000000;
      11'h472: data = 24'b000000000001111100000000;
      11'h473: data = 24'b000000000001111100000000;
      11'h474: data = 24'b000000000001111100000000;
      11'h475: data = 24'b000000000001111100000000;
      11'h476: data = 24'b000000000001111100000000;
      11'h477: data = 24'b000000000001111100000000;
      11'h478: data = 24'b000000000001111100000000;
      11'h479: data = 24'b000000000001111100000000;
      11'h47a: data = 24'b000000000001111100000000;
      11'h47b: data = 24'b000000000001111100000000;
      11'h47c: data = 24'b000000000001111100000000;
      11'h47d: data = 24'b000000000001111100000000;
      11'h47e: data = 24'b000000000001111100000000;
      11'h47f: data = 24'b000000000001111100000000;

      11'h480: data = 24'b000000000000000000000000;
      11'h481: data = 24'b000000000000000000000000;
      11'h482: data = 24'b000000000000000000000000;
      11'h483: data = 24'b000000000000000000000000;
      11'h484: data = 24'b000000000000000000000000;
      11'h485: data = 24'b000000000000000000000000;
      11'h486: data = 24'b000000000000000000000000;
      11'h487: data = 24'b000000000000000000000000;
      11'h488: data = 24'b000000000000000000000000;
      11'h489: data = 24'b000000000000000000000000;
      11'h48a: data = 24'b000000001111111100000000;
      11'h48b: data = 24'b000000111111111111000000;
      11'h48c: data = 24'b000001111111111111110000;
      11'h48d: data = 24'b000011111111111111110000;
      11'h48e: data = 24'b000011111110001111111000;
      11'h48f: data = 24'b000111111000000111111000;
      11'h490: data = 24'b000111110000000011111100;
      11'h491: data = 24'b000111110000000001111100;
      11'h492: data = 24'b001111100000000001111100;
      11'h493: data = 24'b001111100000000001111100;
      11'h494: data = 24'b001111100000000001111100;
      11'h495: data = 24'b000000000000000001111100;
      11'h496: data = 24'b000000000000000001111100;
      11'h497: data = 24'b000000000000000001111100;
      11'h498: data = 24'b000000000000000011111100;
      11'h499: data = 24'b000000000000000011111100;
      11'h49a: data = 24'b000000000000000111111000;
      11'h49b: data = 24'b000000000000000111111000;
      11'h49c: data = 24'b000000000000001111110000;
      11'h49d: data = 24'b000000000000011111110000;
      11'h49e: data = 24'b000000000000011111100000;
      11'h49f: data = 24'b000000000000111111000000;
      11'h4a0: data = 24'b000000000001111110000000;
      11'h4a1: data = 24'b000000000011111110000000;
      11'h4a2: data = 24'b000000000111111100000000;
      11'h4a3: data = 24'b000000001111111000000000;
      11'h4a4: data = 24'b000000011111110000000000;
      11'h4a5: data = 24'b000000111111100000000000;
      11'h4a6: data = 24'b000001111111000000000000;
      11'h4a7: data = 24'b000001111110000000000000;
      11'h4a8: data = 24'b000011111100000000000000;
      11'h4a9: data = 24'b000111111100000000000000;
      11'h4aa: data = 24'b000111111000000000000000;
      11'h4ab: data = 24'b001111110000000000000000;
      11'h4ac: data = 24'b001111111111111111111100;
      11'h4ad: data = 24'b001111111111111111111100;
      11'h4ae: data = 24'b001111111111111111111100;
      11'h4af: data = 24'b011111111111111111111100;

      11'h4b0: data = 24'b000000000000000000000000;
      11'h4b1: data = 24'b000000000000000000000000;
      11'h4b2: data = 24'b000000000000000000000000;
      11'h4b3: data = 24'b000000000000000000000000;
      11'h4b4: data = 24'b000000000000000000000000;
      11'h4b5: data = 24'b000000000000000000000000;
      11'h4b6: data = 24'b000000000000000000000000;
      11'h4b7: data = 24'b000000011111111100000000;
      11'h4b8: data = 24'b000001111111111110000000;
      11'h4b9: data = 24'b000001111111111110000000;
      11'h4ba: data = 24'b000011111111111111000000;
      11'h4bb: data = 24'b000011111000011111110000;
      11'h4bc: data = 24'b001111110000000111110000;
      11'h4bd: data = 24'b001111100000000111111000;
      11'h4be: data = 24'b001111100000000111111000;
      11'h4bf: data = 24'b001111100000000011111000;
      11'h4c0: data = 24'b011111100000000011111000;
      11'h4c1: data = 24'b000000000000000011111000;
      11'h4c2: data = 24'b000000000000000011111000;
      11'h4c3: data = 24'b000000000000000011111000;
      11'h4c4: data = 24'b000000000000000011111000;
      11'h4c5: data = 24'b000000000000000111111000;
      11'h4c6: data = 24'b000000000000001111110000;
      11'h4c7: data = 24'b000000000000011111110000;
      11'h4c8: data = 24'b000000000111111111000000;
      11'h4c9: data = 24'b000000001111111110000000;
      11'h4ca: data = 24'b000000001111111111000000;
      11'h4cb: data = 24'b000000001111111111110000;
      11'h4cc: data = 24'b000000000000001111111000;
      11'h4cd: data = 24'b000000000000000111111100;
      11'h4ce: data = 24'b000000000000000011111100;
      11'h4cf: data = 24'b000000000000000001111100;
      11'h4d0: data = 24'b000000000000000001111110;
      11'h4d1: data = 24'b000000000000000001111110;
      11'h4d2: data = 24'b000000000000000001111110;
      11'h4d3: data = 24'b000000000000000001111110;
      11'h4d4: data = 24'b000000000000000001111110;
      11'h4d5: data = 24'b011111000000000001111110;
      11'h4d6: data = 24'b011111000000000001111110;
      11'h4d7: data = 24'b011111000000000001111100;
      11'h4d8: data = 24'b011111100000000011111100;
      11'h4d9: data = 24'b001111100000000011111100;
      11'h4da: data = 24'b001111110000000111111000;
      11'h4db: data = 24'b000011111000011111111000;
      11'h4dc: data = 24'b000011111111111111110000;
      11'h4dd: data = 24'b000001111111111111000000;
      11'h4de: data = 24'b000001111111111110000000;
      11'h4df: data = 24'b000000011111111100000000;

      11'h4e0: data = 24'b000000000000000000000000;
      11'h4e1: data = 24'b000000000000000000000000;
      11'h4e2: data = 24'b000000000000000000000000;
      11'h4e3: data = 24'b000000000000000000000000;
      11'h4e4: data = 24'b000000000000000000000000;
      11'h4e5: data = 24'b000000000000000000000000;
      11'h4e6: data = 24'b000000000000000000000000;
      11'h4e7: data = 24'b000000000000000000000000;
      11'h4e8: data = 24'b000000000000000000000000;
      11'h4e9: data = 24'b000000000000000000000000;
      11'h4ea: data = 24'b000000000000001111100000;
      11'h4eb: data = 24'b000000000000011111100000;
      11'h4ec: data = 24'b000000000000011111100000;
      11'h4ed: data = 24'b000000000000111111100000;
      11'h4ee: data = 24'b000000000000111111100000;
      11'h4ef: data = 24'b000000000001111111100000;
      11'h4f0: data = 24'b000000000001111111100000;
      11'h4f1: data = 24'b000000000011111111100000;
      11'h4f2: data = 24'b000000000011111111100000;
      11'h4f3: data = 24'b000000000111111111100000;
      11'h4f4: data = 24'b000000001111101111100000;
      11'h4f5: data = 24'b000000001111101111100000;
      11'h4f6: data = 24'b000000011111001111100000;
      11'h4f7: data = 24'b000000011111001111100000;
      11'h4f8: data = 24'b000000111110001111100000;
      11'h4f9: data = 24'b000000111110001111100000;
      11'h4fa: data = 24'b000001111100001111100000;
      11'h4fb: data = 24'b000001111100001111100000;
      11'h4fc: data = 24'b000011111000001111100000;
      11'h4fd: data = 24'b000011111000001111100000;
      11'h4fe: data = 24'b000111110000001111100000;
      11'h4ff: data = 24'b001111100000001111100000;
      11'h500: data = 24'b001111100000001111100000;
      11'h501: data = 24'b011111000000001111100000;
      11'h502: data = 24'b011111000000001111100000;
      11'h503: data = 24'b011111111111111111111110;
      11'h504: data = 24'b011111111111111111111110;
      11'h505: data = 24'b011111111111111111111110;
      11'h506: data = 24'b011111111111111111111110;
      11'h507: data = 24'b000000000000001111100000;
      11'h508: data = 24'b000000000000001111100000;
      11'h509: data = 24'b000000000000001111100000;
      11'h50a: data = 24'b000000000000001111100000;
      11'h50b: data = 24'b000000000000001111100000;
      11'h50c: data = 24'b000000000000001111100000;
      11'h50d: data = 24'b000000000000001111100000;
      11'h50e: data = 24'b000000000000001111100000;
      11'h50f: data = 24'b000000000000001111100000;

      11'h510: data = 24'b000000000000000000000000;
      11'h511: data = 24'b000000000000000000000000;
      11'h512: data = 24'b000000000000000000000000;
      11'h513: data = 24'b000000000000000000000000;
      11'h514: data = 24'b000000000000000000000000;
      11'h515: data = 24'b000000000000000000000000;
      11'h516: data = 24'b000000000000000000000000;
      11'h517: data = 24'b000000000000000000000000;
      11'h518: data = 24'b000000000000000000000000;
      11'h519: data = 24'b000000000000000000000000;
      11'h51a: data = 24'b000000000000000000000000;
      11'h51b: data = 24'b000011111111111111111000;
      11'h51c: data = 24'b000011111111111111111000;
      11'h51d: data = 24'b000011111111111111111000;
      11'h51e: data = 24'b000011111111111111111000;
      11'h51f: data = 24'b000011111000000000000000;
      11'h520: data = 24'b000011111000000000000000;
      11'h521: data = 24'b000111110000000000000000;
      11'h522: data = 24'b000111110000000000000000;
      11'h523: data = 24'b000111110000000000000000;
      11'h524: data = 24'b000111110000000000000000;
      11'h525: data = 24'b000111110000000000000000;
      11'h526: data = 24'b000111110000000000000000;
      11'h527: data = 24'b001111100111111100000000;
      11'h528: data = 24'b001111111111111110000000;
      11'h529: data = 24'b001111111111111111100000;
      11'h52a: data = 24'b001111111111111111110000;
      11'h52b: data = 24'b001111111000011111110000;
      11'h52c: data = 24'b001111110000001111111000;
      11'h52d: data = 24'b001111100000000111111000;
      11'h52e: data = 24'b000000000000000011111000;
      11'h52f: data = 24'b000000000000000011111100;
      11'h530: data = 24'b000000000000000011111100;
      11'h531: data = 24'b000000000000000001111100;
      11'h532: data = 24'b000000000000000001111100;
      11'h533: data = 24'b000000000000000001111100;
      11'h534: data = 24'b000000000000000001111100;
      11'h535: data = 24'b000000000000000011111100;
      11'h536: data = 24'b011111000000000011111100;
      11'h537: data = 24'b011111000000000011111000;
      11'h538: data = 24'b011111100000000011111000;
      11'h539: data = 24'b001111100000000111111000;
      11'h53a: data = 24'b001111110000001111110000;
      11'h53b: data = 24'b001111111100011111110000;
      11'h53c: data = 24'b000111111111111111100000;
      11'h53d: data = 24'b000011111111111111000000;
      11'h53e: data = 24'b000001111111111110000000;
      11'h53f: data = 24'b000000011111111000000000;

      11'h540: data = 24'b000000000000000000000000;
      11'h541: data = 24'b000000000000000000000000;
      11'h542: data = 24'b000000000000000000000000;
      11'h543: data = 24'b000000000000000000000000;
      11'h544: data = 24'b000000000000000000000000;
      11'h545: data = 24'b000000000000000000000000;
      11'h546: data = 24'b000000000000000000000000;
      11'h547: data = 24'b000000000000000000000000;
      11'h548: data = 24'b000000000000000000000000;
      11'h549: data = 24'b000000001111111100000000;
      11'h54a: data = 24'b000000011111111111000000;
      11'h54b: data = 24'b000001111111111111100000;
      11'h54c: data = 24'b000001111111111111100000;
      11'h54d: data = 24'b000011111110011111110000;
      11'h54e: data = 24'b000111111000000111110000;
      11'h54f: data = 24'b000111110000000111111000;
      11'h550: data = 24'b001111110000000011111000;
      11'h551: data = 24'b001111100000000011111000;
      11'h552: data = 24'b001111100000000000000000;
      11'h553: data = 24'b001111100000000000000000;
      11'h554: data = 24'b011111100000000000000000;
      11'h555: data = 24'b011111000000000000000000;
      11'h556: data = 24'b011111000000000000000000;
      11'h557: data = 24'b011111000111111100000000;
      11'h558: data = 24'b011111011111111110000000;
      11'h559: data = 24'b011111111111111111000000;
      11'h55a: data = 24'b011111111111111111100000;
      11'h55b: data = 24'b011111111100011111110000;
      11'h55c: data = 24'b011111111000001111110000;
      11'h55d: data = 24'b011111110000000111111000;
      11'h55e: data = 24'b011111100000000011111000;
      11'h55f: data = 24'b011111100000000011111000;
      11'h560: data = 24'b011111100000000011111100;
      11'h561: data = 24'b011111100000000011111100;
      11'h562: data = 24'b011111000000000001111100;
      11'h563: data = 24'b011111000000000001111100;
      11'h564: data = 24'b011111100000000001111100;
      11'h565: data = 24'b011111100000000011111100;
      11'h566: data = 24'b001111100000000011111100;
      11'h567: data = 24'b001111100000000011111000;
      11'h568: data = 24'b001111110000000011111000;
      11'h569: data = 24'b001111110000000111111000;
      11'h56a: data = 24'b000111111000001111110000;
      11'h56b: data = 24'b000111111110011111110000;
      11'h56c: data = 24'b000011111111111111100000;
      11'h56d: data = 24'b000001111111111111000000;
      11'h56e: data = 24'b000000111111111110000000;
      11'h56f: data = 24'b000000001111111000000000;

      11'h570: data = 24'b000000000000000000000000;
      11'h571: data = 24'b000000000000000000000000;
      11'h572: data = 24'b000000000000000000000000;
      11'h573: data = 24'b000000000000000000000000;
      11'h574: data = 24'b000000000000000000000000;
      11'h575: data = 24'b000000000000000000000000;
      11'h576: data = 24'b000000000000000000000000;
      11'h577: data = 24'b000000000000000000000000;
      11'h578: data = 24'b000000000000000000000000;
      11'h579: data = 24'b000000000000000000000000;
      11'h57a: data = 24'b000000000000000000000000;
      11'h57b: data = 24'b000000000000000000000000;
      11'h57c: data = 24'b011111111111111111111100;
      11'h57d: data = 24'b011111111111111111111100;
      11'h57e: data = 24'b011111111111111111111100;
      11'h57f: data = 24'b011111111111111111111100;
      11'h580: data = 24'b000000000000000111111000;
      11'h581: data = 24'b000000000000000111110000;
      11'h582: data = 24'b000000000000001111110000;
      11'h583: data = 24'b000000000000011111100000;
      11'h584: data = 24'b000000000000011111000000;
      11'h585: data = 24'b000000000000111111000000;
      11'h586: data = 24'b000000000000111110000000;
      11'h587: data = 24'b000000000001111110000000;
      11'h588: data = 24'b000000000001111100000000;
      11'h589: data = 24'b000000000011111100000000;
      11'h58a: data = 24'b000000000011111100000000;
      11'h58b: data = 24'b000000000011111000000000;
      11'h58c: data = 24'b000000000111111000000000;
      11'h58d: data = 24'b000000000111110000000000;
      11'h58e: data = 24'b000000001111110000000000;
      11'h58f: data = 24'b000000001111110000000000;
      11'h590: data = 24'b000000001111100000000000;
      11'h591: data = 24'b000000001111100000000000;
      11'h592: data = 24'b000000011111100000000000;
      11'h593: data = 24'b000000011111000000000000;
      11'h594: data = 24'b000000011111000000000000;
      11'h595: data = 24'b000000011111000000000000;
      11'h596: data = 24'b000000111111000000000000;
      11'h597: data = 24'b000000111110000000000000;
      11'h598: data = 24'b000000111110000000000000;
      11'h599: data = 24'b000000111110000000000000;
      11'h59a: data = 24'b000000111110000000000000;
      11'h59b: data = 24'b000001111110000000000000;
      11'h59c: data = 24'b000001111110000000000000;
      11'h59d: data = 24'b000001111110000000000000;
      11'h59e: data = 24'b000001111100000000000000;
      11'h59f: data = 24'b000001111100000000000000;

      11'h5a0: data = 24'b000000000000000000000000;
      11'h5a1: data = 24'b000000000000000000000000;
      11'h5a2: data = 24'b000000000000000000000000;
      11'h5a3: data = 24'b000000000000000000000000;
      11'h5a4: data = 24'b000000000000000000000000;
      11'h5a5: data = 24'b000000000000000000000000;
      11'h5a6: data = 24'b000000000000000000000000;
      11'h5a7: data = 24'b000000000000000000000000;
      11'h5a8: data = 24'b000000000000000000000000;
      11'h5a9: data = 24'b000000001111111000000000;
      11'h5aa: data = 24'b000000111111111110000000;
      11'h5ab: data = 24'b000001111111111111000000;
      11'h5ac: data = 24'b000011111111111111100000;
      11'h5ad: data = 24'b000111111100011111100000;
      11'h5ae: data = 24'b000111111000001111110000;
      11'h5af: data = 24'b000111110000001111110000;
      11'h5b0: data = 24'b001111110000000111110000;
      11'h5b1: data = 24'b001111100000000111110000;
      11'h5b2: data = 24'b001111100000000111111000;
      11'h5b3: data = 24'b001111100000000111111000;
      11'h5b4: data = 24'b001111100000000111110000;
      11'h5b5: data = 24'b001111110000000111110000;
      11'h5b6: data = 24'b000111110000000111110000;
      11'h5b7: data = 24'b000111111000001111110000;
      11'h5b8: data = 24'b000011111100011111100000;
      11'h5b9: data = 24'b000001111111111111000000;
      11'h5ba: data = 24'b000000111111111110000000;
      11'h5bb: data = 24'b000001111111111110000000;
      11'h5bc: data = 24'b000011111111111111100000;
      11'h5bd: data = 24'b000111111100011111110000;
      11'h5be: data = 24'b001111110000001111110000;
      11'h5bf: data = 24'b001111100000000111111000;
      11'h5c0: data = 24'b011111100000000011111000;
      11'h5c1: data = 24'b011111000000000011111000;
      11'h5c2: data = 24'b011111000000000011111100;
      11'h5c3: data = 24'b011111000000000001111100;
      11'h5c4: data = 24'b011111000000000001111100;
      11'h5c5: data = 24'b011111000000000001111100;
      11'h5c6: data = 24'b011111000000000011111100;
      11'h5c7: data = 24'b011111100000000011111100;
      11'h5c8: data = 24'b011111100000000011111000;
      11'h5c9: data = 24'b001111110000000111111000;
      11'h5ca: data = 24'b001111110000001111111000;
      11'h5cb: data = 24'b000111111100011111110000;
      11'h5cc: data = 24'b000111111111111111100000;
      11'h5cd: data = 24'b000011111111111111000000;
      11'h5ce: data = 24'b000000111111111110000000;
      11'h5cf: data = 24'b000000001111111000000000;

      11'h5d0: data = 24'b000000000000000000000000;
      11'h5d1: data = 24'b000000000000000000000000;
      11'h5d2: data = 24'b000000000000000000000000;
      11'h5d3: data = 24'b000000000000000000000000;
      11'h5d4: data = 24'b000000000000000000000000;
      11'h5d5: data = 24'b000000000000000000000000;
      11'h5d6: data = 24'b000000000000000000000000;
      11'h5d7: data = 24'b000000000000000000000000;
      11'h5d8: data = 24'b000000000000000000000000;
      11'h5d9: data = 24'b000000011111110000000000;
      11'h5da: data = 24'b000000111111111100000000;
      11'h5db: data = 24'b000011111111111110000000;
      11'h5dc: data = 24'b000011111111111111000000;
      11'h5dd: data = 24'b000111111100011111100000;
      11'h5de: data = 24'b001111111000001111110000;
      11'h5df: data = 24'b001111110000000111110000;
      11'h5e0: data = 24'b001111100000000111110000;
      11'h5e1: data = 24'b011111100000000011111000;
      11'h5e2: data = 24'b011111000000000011111000;
      11'h5e3: data = 24'b011111000000000011111000;
      11'h5e4: data = 24'b011111000000000011111000;
      11'h5e5: data = 24'b011111000000000011111000;
      11'h5e6: data = 24'b011111000000000011111100;
      11'h5e7: data = 24'b011111000000000011111100;
      11'h5e8: data = 24'b011111000000000011111100;
      11'h5e9: data = 24'b011111100000000011111100;
      11'h5ea: data = 24'b011111100000000111111100;
      11'h5eb: data = 24'b001111110000000111111100;
      11'h5ec: data = 24'b001111110000001111111100;
      11'h5ed: data = 24'b000111111100011111111100;
      11'h5ee: data = 24'b000111111111111111111100;
      11'h5ef: data = 24'b000011111111111101111100;
      11'h5f0: data = 24'b000001111111111001111100;
      11'h5f1: data = 24'b000000011111110011111100;
      11'h5f2: data = 24'b000000000000000011111000;
      11'h5f3: data = 24'b000000000000000011111000;
      11'h5f4: data = 24'b000000000000000011111000;
      11'h5f5: data = 24'b000000000000000011111000;
      11'h5f6: data = 24'b000000000000000111111000;
      11'h5f7: data = 24'b001111100000000111110000;
      11'h5f8: data = 24'b001111100000000111110000;
      11'h5f9: data = 24'b001111100000001111110000;
      11'h5fa: data = 24'b001111110000011111100000;
      11'h5fb: data = 24'b000111111000111111100000;
      11'h5fc: data = 24'b000111111111111111000000;
      11'h5fd: data = 24'b000011111111111110000000;
      11'h5fe: data = 24'b000001111111111100000000;
      11'h5ff: data = 24'b000000011111110000000000;
		
		11'h600: data = 24'b000000000000000000000000;
      11'h601: data = 24'b000000000000000000000000;
      11'h602: data = 24'b000000000000000000000000;
      11'h603: data = 24'b000000000000000000000000;
      11'h604: data = 24'b000000000000000000000000;
      11'h605: data = 24'b000000000000000000000000;
      11'h606: data = 24'b000000000000000000000000;
      11'h607: data = 24'b000000000000000000000000;
      11'h608: data = 24'b000000000000000000000000;
      11'h609: data = 24'b000000000000000000000000;
      11'h60a: data = 24'b000000000000000000000000;
      11'h60b: data = 24'b000000000000000000000000;
      11'h60c: data = 24'b000000001111110000000000;
      11'h60d: data = 24'b000000001111110000000000;
      11'h60e: data = 24'b000000001111110000000000;
      11'h60f: data = 24'b000000001111110000000000;
      11'h610: data = 24'b000000001111110000000000;
      11'h611: data = 24'b000000000000000000000000;
      11'h612: data = 24'b000000000000000000000000;
      11'h613: data = 24'b000000000000000000000000;
      11'h614: data = 24'b000000000000000000000000;
      11'h615: data = 24'b000000000000000000000000;
      11'h616: data = 24'b000000000000000000000000;
      11'h617: data = 24'b000000000000000000000000;
      11'h618: data = 24'b000000000000000000000000;
      11'h619: data = 24'b000000000000000000000000;
      11'h61a: data = 24'b000000000000000000000000;
      11'h61b: data = 24'b000000000000000000000000;
      11'h61c: data = 24'b000000000000000000000000;
      11'h61d: data = 24'b000000000000000000000000;
      11'h61e: data = 24'b000000000000000000000000;
      11'h61f: data = 24'b000000000000000000000000;
      11'h620: data = 24'b000000000000000000000000;
      11'h621: data = 24'b000000001111110000000000;
      11'h622: data = 24'b000000001111110000000000;
      11'h623: data = 24'b000000001111110000000000;
      11'h624: data = 24'b000000001111110000000000;
      11'h625: data = 24'b000000001111110000000000;
      11'h626: data = 24'b000000000000000000000000;
      11'h627: data = 24'b000000000000000000000000;
      11'h628: data = 24'b000000000000000000000000;
      11'h629: data = 24'b000000000000000000000000;
      11'h62a: data = 24'b000000000000000000000000;
      11'h62b: data = 24'b000000000000000000000000;
      11'h62c: data = 24'b000000000000000000000000;
      11'h62d: data = 24'b000000000000000000000000;
      11'h62e: data = 24'b000000000000000000000000;
      11'h62f: data = 24'b000000000000000000000000;
		
		11'h630: data = 24'b000000000000000000000000;
      11'h631: data = 24'b000000000000000000000000;
      11'h632: data = 24'b000000000000000000000000;
      11'h633: data = 24'b000000000000000000000000;
      11'h634: data = 24'b000000000000000000000000;
      11'h635: data = 24'b000000000000000000000000;
      11'h636: data = 24'b000000000000000000000000;
      11'h637: data = 24'b000000000000000000000000;
      11'h638: data = 24'b000000000000000000000000;
      11'h639: data = 24'b000000000000000000000000;
      11'h63a: data = 24'b000000000000000000000000;
      11'h63b: data = 24'b000000000000000000000000;
      11'h63c: data = 24'b000000000000000000000000;
      11'h63d: data = 24'b000000000000000000000000;
      11'h63e: data = 24'b000000000000000000000000;
      11'h63f: data = 24'b000000000000000000000000;
      11'h640: data = 24'b000000000000000000000000;
      11'h641: data = 24'b000000000000000000000000;
      11'h642: data = 24'b011111000111110000000000;
      11'h643: data = 24'b111111101111111000000000;
      11'h644: data = 24'b111111111111111000000000;
      11'h645: data = 24'b111111111111111000000000;
      11'h646: data = 24'b111111111111111000000000;
      11'h647: data = 24'b111111111111111000000000;
      11'h648: data = 24'b111111111111110000000000;
      11'h649: data = 24'b011111111111110000000000;
      11'h64a: data = 24'b011111111111100000000000;
      11'h64b: data = 24'b001111111111000000000000;
      11'h64c: data = 24'b000111111110000000000000;
      11'h64d: data = 24'b000011111100000000000000;
      11'h64e: data = 24'b000001111000000000000000;
      11'h64f: data = 24'b000000110000000000000000;
      11'h650: data = 24'b000000000000000000000000;
      11'h651: data = 24'b000000000000000000000000;
      11'h652: data = 24'b000000000000000000000000;
      11'h653: data = 24'b000000000000000000000000;
      11'h654: data = 24'b000000000000000000000000;
      11'h655: data = 24'b000000000000000000000000;
      11'h656: data = 24'b000000000000000000000000;
      11'h657: data = 24'b000000000000000000000000;
      11'h658: data = 24'b000000000000000000000000;
      11'h659: data = 24'b000000000000000000000000;
      11'h65a: data = 24'b000000000000000000000000;
      11'h65b: data = 24'b000000000000000000000000;
      11'h65c: data = 24'b000000000000000000000000;
      11'h65d: data = 24'b000000000000000000000000;
      11'h65e: data = 24'b000000000000000000000000;
      11'h65f: data = 24'b000000000000000000000000;
		
		11'h660: data = 24'b000000000000000000000000;
      11'h661: data = 24'b000000000000000000000000;
      11'h662: data = 24'b000000000000000000000000;
      11'h663: data = 24'b000000000000000000000000;
      11'h664: data = 24'b000000000000000000000000;
      11'h665: data = 24'b000000000000000000000000;
      11'h666: data = 24'b000000000000000000000000;
      11'h667: data = 24'b000000000000000000000000;
      11'h668: data = 24'b000000000000000000000000;
      11'h669: data = 24'b000000000000000000000000;
      11'h66a: data = 24'b000000000001110000000000;
      11'h66b: data = 24'b000000000011110000000000;
      11'h66c: data = 24'b000000000011100000000000;
      11'h66d: data = 24'b000000000011100000000000;
      11'h66e: data = 24'b000000000111100000000000;
      11'h66f: data = 24'b000000000111000000000000;
      11'h670: data = 24'b000000001111000000000000;
      11'h671: data = 24'b000000001110000000000000;
      11'h672: data = 24'b000000011110000000000000;
      11'h673: data = 24'b000000011110000000000000;
      11'h674: data = 24'b000000011100000000000000;
      11'h675: data = 24'b000000111100000000000000;
      11'h676: data = 24'b000000111000000000000000;
      11'h677: data = 24'b000001111000000000000000;
      11'h678: data = 24'b000001111000000000000000;
      11'h679: data = 24'b000001110000000000000000;
      11'h67a: data = 24'b000011110000000000000000;
      11'h67b: data = 24'b000011100000000000000000;
      11'h67c: data = 24'b000111100000000000000000;
      11'h67d: data = 24'b000111000000000000000000;
      11'h67e: data = 24'b001111000000000000000000;
      11'h67f: data = 24'b001111000000000000000000;
      11'h680: data = 24'b000000000000000000000000;
      11'h681: data = 24'b000000000000000000000000;
      11'h682: data = 24'b000000000000000000000000;
      11'h683: data = 24'b000000000000000000000000;
      11'h684: data = 24'b000000000000000000000000;
      11'h685: data = 24'b000000000000000000000000;
      11'h686: data = 24'b000000000000000000000000;
      11'h687: data = 24'b000000000000000000000000;
      11'h688: data = 24'b000000000000000000000000;
      11'h689: data = 24'b000000000000000000000000;
      11'h68a: data = 24'b000000000000000000000000;
      11'h68b: data = 24'b000000000000000000000000;
      11'h68c: data = 24'b000000000000000000000000;
      11'h68d: data = 24'b000000000000000000000000;
      11'h68e: data = 24'b000000000000000000000000;
      11'h68f: data = 24'b000000000000000000000000;
		
		11'h690: data = 24'b000000000000000000000000;
      11'h691: data = 24'b000000000000000000000000;
      11'h692: data = 24'b000000000000000000000000;
      11'h693: data = 24'b000000000000000000000000;
      11'h694: data = 24'b000000000000000000000000;
      11'h695: data = 24'b000000000000000000000000;
      11'h696: data = 24'b000000000000000000000000;
      11'h697: data = 24'b000000000000000000000000;
      11'h698: data = 24'b000000000000000000000000;
      11'h699: data = 24'b000000000000000000000000;
      11'h69a: data = 24'b000000000000000000000000;
      11'h69b: data = 24'b000000000000000000000000;
      11'h69c: data = 24'b011110111111000000000000;
      11'h69d: data = 24'b011111111111110000000000;
      11'h69e: data = 24'b011111100011110000000000;
      11'h69f: data = 24'b011111000001111000000000;
      11'h6a0: data = 24'b011110000001111000000000;
      11'h6a1: data = 24'b011110000000111000000000;
      11'h6a2: data = 24'b011110000000111000000000;
      11'h6a3: data = 24'b011110000000111000000000;
      11'h6a4: data = 24'b011110000000111000000000;
      11'h6a5: data = 24'b011110000001111000000000;
      11'h6a6: data = 24'b011111000001111000000000;
      11'h6a7: data = 24'b011111100011110000000000;
      11'h6a8: data = 24'b011111111111100000000000;
      11'h6a9: data = 24'b011110111111000000000000;
      11'h6aa: data = 24'b011110000000000000000000;
      11'h6ab: data = 24'b011110000000000000000000;
      11'h6ac: data = 24'b011110000000000000000000;
      11'h6ad: data = 24'b011110000000000000000000;
      11'h6ae: data = 24'b011110000000000000000000;
      11'h6af: data = 24'b011110000000000000000000;
      11'h6b0: data = 24'b000000000000000000000000;
      11'h6b1: data = 24'b000000000000000000000000;
      11'h6b2: data = 24'b000000000000000000000000;
      11'h6b3: data = 24'b000000000000000000000000;
      11'h6b4: data = 24'b000000000000000000000000;
      11'h6b5: data = 24'b000000000000000000000000;
      11'h6b6: data = 24'b000000000000000000000000;
      11'h6b7: data = 24'b000000000000000000000000;
      11'h6b8: data = 24'b000000000000000000000000;
      11'h6b9: data = 24'b000000000000000000000000;
      11'h6ba: data = 24'b000000000000000000000000;
      11'h6bb: data = 24'b000000000000000000000000;
      11'h6bc: data = 24'b000000000000000000000000;
      11'h6bd: data = 24'b000000000000000000000000;
      11'h6be: data = 24'b000000000000000000000000;
      11'h6bf: data = 24'b000000000000000000000000;
		
		11'h6c0: data = 24'b000000000000000000000000;
      11'h6c1: data = 24'b000000000000000000000000;
      11'h6c2: data = 24'b000000000000000000000000;
      11'h6c3: data = 24'b000000000000000000000000;
      11'h6c4: data = 24'b000000000000000000000000;
      11'h6c5: data = 24'b000000000000000000000000;
      11'h6c6: data = 24'b000000000000000000000000;
      11'h6c7: data = 24'b000000000000000000000000;
      11'h6c8: data = 24'b000000000000000000000000;
      11'h6c9: data = 24'b000000000000000000000000;
      11'h6ca: data = 24'b000000000000000000000000;
      11'h6cb: data = 24'b000000000000000000000000;
      11'h6cc: data = 24'b000000000000000000000000;
      11'h6cd: data = 24'b000000000000000000000000;
      11'h6ce: data = 24'b000000000000000000000000;
      11'h6cf: data = 24'b000000000000000000000000;
      11'h6d0: data = 24'b000000000000000000000000;
      11'h6d1: data = 24'b000000000000000000000000;
      11'h6d2: data = 24'b000000000000000000000000;
      11'h6d3: data = 24'b000000000000000000000000;
      11'h6d4: data = 24'b000000000000000000000000;
      11'h6d5: data = 24'b000000000000000000000000;
      11'h6d6: data = 24'b000000000000000000000000;
      11'h6d7: data = 24'b000000000000000000000000;
      11'h6d8: data = 24'b000000000000000000000000;
      11'h6d9: data = 24'b000000000000000000000000;
      11'h6da: data = 24'b000000000000000000000000;
      11'h6db: data = 24'b000000000000000000000000;
      11'h6dc: data = 24'b000000000000000000000000;
      11'h6dd: data = 24'b000000000000000000000000;
      11'h6de: data = 24'b000000000000000000000000;
      11'h6df: data = 24'b000000000000000000000000;
      11'h6e0: data = 24'b000000000000000000000000;
      11'h6e1: data = 24'b000000000000000000000000;
      11'h6e2: data = 24'b000000000000000000000000;
      11'h6e3: data = 24'b000000000000000000000000;
      11'h6e4: data = 24'b000000000000000000000000;
      11'h6e5: data = 24'b000000000000000000000000;
      11'h6e6: data = 24'b000000000000000000000000;
      11'h6e7: data = 24'b000000000000000000000000;
      11'h6e8: data = 24'b000000000000000000000000;
      11'h6e9: data = 24'b000000000000000000000000;
      11'h6ea: data = 24'b000000000000000000000000;
      11'h6eb: data = 24'b000000000000000000000000;
      11'h6ec: data = 24'b000000000000000000000000;
      11'h6ed: data = 24'b000000000000000000000000;
      11'h6ee: data = 24'b000000000000000000000000;
      11'h6ef: data = 24'b000000000000000000000000;






    endcase
end

endmodule
